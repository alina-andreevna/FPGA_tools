----------------------------------------------------------------------------------
-- MOD.DATE: 
--------------------------------------------------
-- Project :		
-- Author :			Alina Galichina
-- Creation date : 	
-- File : 			.vhd
-- TestBench : 		..\_tb.vhd
-- Software : 		ISE 14.7, Vivado 2018
-- Primitives : 	No
-- Cores : 			No
-- Submodules : 	No
--------------------------------------------------
-- Description : 	
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity <entity_name> is

	generic(
		);    

	port( clk        : in  std_logic;
		  rst_in     : in std_logic;

		  _in			: in std_logic;
		  _in			: in std_logic_vector( downto );

		  _out			: out std_logic;
		  _out			: out std_logic_vector( downto );	

		  );

end entity <entity_name>;

--------------------------------------------------

architecture <arch_name> of <entity_name> is

	------------------=FUNCTIONS=------------------

-- NO FUCTIONS --

	------------------=END FUNCTIONS=------------------


	------------------=CONSTANTS,SIGNALS,VARIABLES=------------------

-- NO SIGNALS, CONSTANTS AND VARIABLES --
	
	------------------=END CONSTANTS,SIGNALS,VARIABLES=------------------


	-----------------=COMPONENTS=------------------

-- NO COMPONENTS --

	------------------=END COMPONENTS=------------------


	-----------------=DEBUG ZONE=------------------

-- NO DEBUG ZONE --

	------------------=END DEBUG ZONE=------------------


	-----------------=ATTRIBUTES=------------------

-- NO ATTRIBUTES --

	------------------=END ATTRIBUTES=------------------

--------------------------------------------------

begin

	----=ASSERTIONS=----

-- NO ASSERTIONS --

	----=END ASSERTIONS=----


	----=CONTINIOUS ASSIGNMENTS=----

-- NO CONTINIOUS ASSIGNMENTS --

	----=END CONTINIOUS ASSIGNMENTS=----


	----=INSTANCES=---

-- NO INSTANCES --

	----=END INSTANCES=----


	----=PROCESSES ETC.=----
	
-- NO PROCESSES ETC. --

	----=END PROCESSES ETC.=----


	----=DEBUG ZONE=----

-- NO DEBUG ZONE --

	----=END DEBUG ZONE=----

end architecture <arch_name>;